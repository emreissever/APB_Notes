`timescale 1ns / 1ps

module APB_MasterModule_Tb();

reg clk = 1;
reg rstN = 1; 

reg [31:0]      apb_addr;
reg             apb_write;
reg             apb_sel;
reg             apb_en;
reg [31:0]      apb_wdata;

wire            apb_rdata;
wire            apb_ready;
wire            pwm_out;


APB_PWM APB_PWM_Test
(
    .PCLK(clk),
    .PRESETn(rstN),

    .PADDR(apb_addr),
    .PWRITE(apb_write),
    .PSEL(apb_sel),
    .PENABLE(apb_en),
    .PWDATA(apb_wdata),

    .PREADY(apb_ready),

    .PWM_OUT(pwm_out)
);

always
// CLOCK Period = 62.5 ns 
// Assumed Controller Frequency Is 16 MHz (Arduino)
#(31.25) clk = !clk;
initial begin

    // Initial values
    clk = 1;
    rstN = 1;
    apb_sel   = 0;
    apb_en    = 0;
    apb_addr  = 0;
    apb_wdata  = 0;
    apb_write = 0;
/* 
    // First Write
    @(posedge clk);
    apb_sel   = 1;
    apb_write = 1;
    apb_addr  = 1;
    apb_wdata  = 120;
    @(posedge clk);
    apb_en = 1;
    @(posedge clk); 
    if(apb_ready) begin
        apb_en    = 0;
        apb_addr  = 2;
        apb_wdata  = 5;
    end
    else begin
        $display("Timeout"); 
    end

    // Second Write
    @(posedge clk);
    apb_en = 1;
    @(posedge clk); 
    if(apb_ready) begin
        apb_en    = 0;
        apb_sel   = 1;
        apb_addr  = 0;
        apb_wdata  = 1;
    end

    @(posedge clk);
    apb_en = 1;
    @(posedge clk); 
    if(apb_ready) begin
        apb_en    = 0;
        apb_sel   = 0;
        apb_addr  = 0;
        apb_wdata  = 0;
        $display("Success");
    end
    else begin
        $display("Failed TimeOut");
    end
 */
/*     @(posedge clk);
    apb_en    = 0;
    apb_sel   = 0; */
    #625;
    //#2000;
    $finish;
end

// 'Memory Address', 'Write Data' and 'Multiple Write' as Input 
task write_transfer(input [31:0] MemAddr, input [31:0] WriteData, input mulWrite);
begin
    @(posedge clk);
    apb_sel    = 1;
    apb_write  = 1;
    apb_addr   = MemAddr;
    apb_wdata  = WriteData;
    @(posedge clk);
    apb_en = 1;
    @(posedge clk);
    if(apb_ready) begin
        apb_en = 0; 
        if(~mulWrite) apb_sel = 0;
    end
end
endtask
endmodule
